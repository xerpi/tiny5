package cache_interface_types;

typedef enum logic [1:0] {
	CACHE_ACCESS_SIZE_BYTE,
	CACHE_ACCESS_SIZE_HALF,
	CACHE_ACCESS_SIZE_WORD
} cache_access_size_t;

endpackage
